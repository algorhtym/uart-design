library ieee;
use ieee.std_logic_1164.all;

entity tx_control is
    port (
   
    );
end tx_control;

-- FSM :
--      s1 --[]


architecture struc_tx_control of tx_control is

    -- signal declarations

    -- component declarations



begin
    -- components

    -- signal connections

    -- output driver
    

end struc_tx_control;