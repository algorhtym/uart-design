library ieee;
use ieee.std_logic_1164.all;

entity transmitter_control is
    port (
        reset_bar : in std_logic;


    );

    -- s1 : 